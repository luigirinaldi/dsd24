module cordic_cos #(
    parameter NUM_ITER = 20,
    parameter FRAC_BITS = 20
)

(
    input signed wire [FRAC_BITS+1:0] theta_in,
    output signed wire [FRAC_BITS+1:0] cos_out
)



endmodule